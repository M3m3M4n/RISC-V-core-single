/* Flag behaviours:  http://personal.denison.edu/~bressoud/cs281-s08/homework/MIPSALU.html
 * Comparison:       https://people.cs.pitt.edu/~don/coe1502/current/Unit1/CompBlock/ALU_Comp.html
 * Overflow / carry: http://teaching.idallen.com/dat2343/10f/notes/040_overflow.txt
 * Subtract / comp:  https://mil.ufl.edu/3701/classes/11%20Add,%20Subtract,%20Compare,%20ALU.pdf
 */

module ALU (
    input  logic [31:0] a, b,
    input  logic [3:0]  alu_control,
    output logic [31:0] result,
    output logic [3:0]  alu_flags
);

    logic zero;
    logic neg;
    logic carry;
    logic overflow;

    logic [31:0] condinvb;
    logic [32:0] sum;
    logic        isAddSub; // true when is add or subtract operation
    logic        isSub;

    assign alu_flags[0] = zero;
    assign alu_flags[1] = neg;
    assign alu_flags[2] = carry;
    assign alu_flags[3] = overflow;

    /* Condition for subtraction must also statisfy when slt and sltu is active
     * Range from 4'b0000 to 4'b0011
     */
    assign isAddSub = ~alu_control[2] & ~alu_control[3];
    assign isSub    = isAddSub & (alu_control[0] | alu_control[1]);
    assign condinvb = isSub ? ~b : b;
    
    assign sum      = a + condinvb + isSub;

    assign zero     = (result == 32'b0);
    assign neg      = (result[31] == 1'b1);
    assign overflow = ~(isSub ^ a[31] ^ b[31]) & (a[31] ^ sum[31]) & isAddSub;

    /* Assumption about subtraction carry (borrow)
     * If addition of 2's complement result in carry => no subtraction carry
     * Else if addition does not result in a carry => subtraction carry
     * Boolean: isSub = C; sum[32] = S
     * Need prove: (C & ~S) | (~C & S) => C^S
     * Consider adding 2 complement = adding inverse bit with initial carry = 1
     * Subtraction: B(i+1) = ~MiSi + ~MiBi + SiBi
     * Add 2 complement: C(i+1) = Mi~Si + MiCi + ~SiCi
     * Assumption: B(out) == ~C(out)
     * ~C(i+1) = ~MiSi + ~Mi~Ci + Si~Ci => maybe prove by recursive back to C0 = 1 vs B0 = 0?
     */
    assign carry    = (isSub ^ sum[32]) & isAddSub;

    always_comb begin
        case (alu_control)
            4'b0000: result = sum[31:0];          // add
            4'b0001: result = sum[31:0];          // subtract
            4'b0010: result = sum[31] ^ overflow; // slt
            4'b0011: result = carry;              // sltu
            4'b0100: result = a ^ b;              // xor
            4'b0101: result = a & b;              // and 
            4'b0110: result = a | b;              // or
            4'b0111: result = a << b[4:0];        // sll
            4'b1000: result = a >> b[4:0];        // srl
            4'b1001: result = a >>> b[4:0];       // sra
            default: result = 32'bx;
        endcase
    end

endmodule